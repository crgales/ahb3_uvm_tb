package ahb_env_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import ahb_agent_pkg::*;
  `include "ahb_env_config.svh"
  `include "ahb_coverage.svh"
  `include "ahb_env.svh"
endpackage