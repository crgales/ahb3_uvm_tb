package ahb_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import ahb_agent_pkg::*;
  import ahb_env_pkg::*;

  `include "ahb_base_vseq.svh"
  `include "ahb_vseq.svh"
  `include "ahb_base_test.svh"
  `include "ahb_simple_test.svh"
endpackage